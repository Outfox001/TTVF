// ------------------------------------------------------------------------------------------------------------------------------------------------------------------------
// Module name: afvip_test_pkg
// HDL        : UVM
// Author     : Paulovici Vlad-Marian
// Description: Package for the library of tests and virtual sequence
// Date       : 28 August, 2023
// -----------------------------------------------------------------------------------------------------------------------------------------------------------------------------


package test_pkg;

  import uvm_pkg::*;
  import apb_pkg::*;
  import reset_pkg::*;
  import output_pkg::*;
  import env_pkg::*;

  `include "uvm_macros.svh"
  `include "test_lib.svh"
   
endpackage