// ------------------------------------------------------------------------------------------------------------------------------------------------------------------------
// Module name: reset_pkg
// HDL        : System Verilog
// Author     : Paulovici Vlad-Marian
// Description: Package for reset
// Date       : 28 August, 2023
// -----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
package reset_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "reset_item.svh"
  `include "reset_driver.svh"
  `include "reset_monitor.svh"
  `include "reset_sequencer.svh"
  `include "reset_agent.svh"
  `include "reset_sequence.svh"
    
endpackage